library verilog;
use verilog.vl_types.all;
entity decoder_2_4_vlg_vec_tst is
end decoder_2_4_vlg_vec_tst;
